** Profile: "SCHEMATIC1-myfinalsimu"  [ c:\analog circuits assigments\updated_project\finalupdatedproject-PSpiceFiles\SCHEMATIC1\myfinalsimu.sim ] 

** Creating circuit file "myfinalsimu.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../finalupdatedproject-pspicefiles/finalupdatedproject.lib" 
* From [PSPICE NETLIST] section of C:\Users\orsha\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100000 100 110000000
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
